`include "define.v"
module rom (
    input addr_i,
    input ce,
    output addr_o,
    output inst
);
    
    
endmodule
`include "buceros_header.v"
module ram (
    input [`InstAddrBus] addr,
    input we,
    input re,
    input sel,
    input data_i,
    input ce,
    input rst,
    input clk,
    output data_o
);

    
endmodule
/*
 * Description  : Bus Interface Unit
 * Author       : Zhengyi Zhang
 * Date         : 2021-11-25 17:10:47
 * LastEditTime : 2021-11-28 13:16:30
 * LastEditors  : Zhengyi Zhang
 * FilePath     : \Buceros\src\core\biu.v
 */
module biu (
);

endmodule //biu
module rom (
    input  wire                clk,
);
    
endmodule
module uart_top (
);

endmodule //uart_top